module debug_rom(
    input wire clk,
    input wire rstn,
    input wire[31:0] addr,
    input wire addr_valid,
    output wire addr_ready,
    output reg rvalid,
    output reg[31:0] rdata
);

    wire[31:0] rom_content[22] = '{
        32'h7b241073, // csrw dscratch0, s0
        32'h10002023, // sw x0, HALTED
        32'h10806403, // lwu s0, GOING
        32'h04041063, // bnez s0S, 64
        32'h11006403, // lwu s0, ACK
        32'hfe040ae3, // beqz s0, -12

        32'h10002823, // sw x0, ACK
        32'h7b349073, // csrw dscratch1, s1
        32'h00100413, // li s0, 1
        32'h01441493, // li s1, 0x0010_0000
        32'h01f41413, // li s0, 0x8000_0000
        32'h009464b3, // li s1, 0x8010_0000
        32'h00040003, // lb x0, 0(s0)
        32'h01040413, // addi	s0,s0,16
        32'hfe941ce3, // bne	s0,s1,-8
        32'h7b3024f3, // csrr s1, dscratch1
        32'h7b206473, // csrr s0, dscratch0
        32'h10002c23, // sw x0, RESUME
        32'h7b200073, // dret

        32'h7b206473, // csrr s0, dscratch0
        32'h10002423, // sw x0, GOING
        32'h30000067  // j 0x300 jumps to abstract command
    };
    always_ff @(posedge clk or negedge rstn)
        if (!rstn)
            rvalid <= 1'b0;
        else
            rvalid <= addr_valid & addr_ready;

    always_ff @(posedge clk or negedge rstn)
        if (!rstn)
            rdata <= '0;
        else if (addr_valid & addr_ready)
            rdata <= rom_content[addr[31:2]];
    
    assign addr_ready = 1'b1;
    

endmodule


module boot_rom(
    input wire clk,
    input wire rstn,
    input wire[31:0] addr,
    input wire addr_valid,
    output wire addr_ready,
    output reg rvalid,
    output reg[31:0] rdata,

    input wire[31:0] addr2,
    input wire addr2_valid,
    output wire addr2_ready,
    output reg rvalid2,
    output reg[63:0] rdata2
    
);

    wire[31:0] rom_content[335] = '{32'h70001137,
32'h70000437,
32'h700014b7,
32'h00843023,
32'h00840413,
32'hfe941ce3,
32'h70000437,
32'h00043503,
32'h00851c63,
32'h00840413,
32'hfe941ae3,
32'h010000ef,
32'h700000b7,
32'h00008067,
32'h0000006f,
32'hfb010113,
32'h00000517,
32'h48050513,
32'h04813023,
32'h02913c23,
32'h04113423,
32'h03213823,
32'h03313423,
32'h03413023,
32'h01513c23,
32'h37c000ef,
32'h100247b7,
32'h0a600713,
32'h00e7a023,
32'h01878413,
32'h00300793,
32'h00f42023,
32'h00a00493,
32'hfff48493,
32'h2dc000ef,
32'hfe049ce3,
32'h00000517,
32'h44050513,
32'h00042023,
32'h344000ef,
32'h09500613,
32'h00000593,
32'h04000513,
32'h358000ef,
32'h00050913,
32'h2b8000ef,
32'h00100793,
32'h26f91863,
32'h00000517,
32'h41850513,
32'h318000ef,
32'h08700613,
32'h1aa00593,
32'h04800513,
32'h32c000ef,
32'h0005049b,
32'h284000ef,
32'h280000ef,
32'h27c000ef,
32'h00050413,
32'h274000ef,
32'h0005051b,
32'hfff48493,
32'hf5650513,
32'h00f47413,
32'h009034b3,
32'h00a03533,
32'hfff40413,
32'h00a4e4b3,
32'h00803433,
32'h00946433,
32'h250000ef,
32'h20041663,
32'h00000517,
32'h3bc50513,
32'h2b4000ef,
32'h06500613,
32'h00000593,
32'h07700513,
32'h2c8000ef,
32'h22c000ef,
32'h07700613,
32'h400005b7,
32'h06900513,
32'h2b4000ef,
32'hfd250ee3,
32'h1c051a63,
32'h00000517,
32'h38c50513,
32'h27c000ef,
32'h0fd00613,
32'h00000593,
32'h07a00513,
32'h290000ef,
32'h00050413,
32'h1e8000ef,
32'hfff54793,
32'h0ff7f793,
32'h0077d79b,
32'h00803433,
32'h00f46433,
32'h1d0000ef,
32'h1cc000ef,
32'h1c8000ef,
32'h1cc000ef,
32'h18041463,
32'h00000517,
32'h34850513,
32'h230000ef,
32'h01500613,
32'h20000593,
32'h05000513,
32'h244000ef,
32'h00a13423,
32'h1a4000ef,
32'h00813503,
32'h14051e63,
32'h00000517,
32'h32450513,
32'h204000ef,
32'h00000517,
32'h32050513,
32'h1c4000ef,
32'h100247b7,
32'h00300713,
32'h00e7a023,
32'h0e100613,
32'h00000593,
32'h05200513,
32'h200000ef,
32'h700009b7,
32'h10051e63,
32'h000024b7,
32'h70001437,
32'h0fe00913,
32'hfe048493,
32'hc0040413,
32'h140000ef,
32'hff251ee3,
32'h00000a13,
32'h20098a93,
32'h130000ef,
32'h00098793,
32'h00a78023,
32'h008a579b,
32'h008a1a1b,
32'h014787b3,
32'h00f547b3,
32'h03079793,
32'h0307d793,
32'h0047d71b,
32'h00f77713,
32'h00e7c7b3,
32'h0107979b,
32'h4107d79b,
32'h00c7971b,
32'h00e7c7b3,
32'h0107979b,
32'h4107d79b,
32'h0057971b,
32'h00977733,
32'h00e7c7b3,
32'h03079a13,
32'h00198993,
32'h030a5a13,
32'hfb5990e3,
32'h0cc000ef,
32'h02851793,
32'h4287da93,
32'h008a9a93,
32'h0bc000ef,
32'h01556533,
32'h03051513,
32'h03055513,
32'h09450263,
32'h00000517,
32'h25450513,
32'h11c000ef,
32'h00100413,
32'h0a0000ef,
32'h00100613,
32'h00000593,
32'h04c00513,
32'h128000ef,
32'h08c000ef,
32'h00000517,
32'h24450513,
32'h0f4000ef,
32'h02041e63,
32'h00000517,
32'h24450513,
32'h0e4000ef,
32'h04813083,
32'h04013403,
32'h03813483,
32'h03013903,
32'h02813983,
32'h02013a03,
32'h01813a83,
32'h00000513,
32'h05010113,
32'h00008067,
32'h044000ef,
32'h00000517,
32'h20450513,
32'h0ac000ef,
32'h0000006f,
32'hee8994e3,
32'h00000413,
32'hf89ff06f,
32'h100247b7,
32'h04a7a423,
32'h04c78793,
32'h0007a703,
32'hfe074ee3,
32'h0ff77513,
32'h00008067,
32'h0ff00513,
32'hfe1ff06f,
32'hff010113,
32'h00113423,
32'hff1ff0ef,
32'h00813083,
32'h100247b7,
32'h0007ac23,
32'h01010113,
32'h00008067,
32'h100137b7,
32'h00100713,
32'h00e7a423,
32'h0007a703,
32'hfe071ee3,
32'h0005051b,
32'h00a7a023,
32'h00008067,
32'hff010113,
32'h00813023,
32'h00113423,
32'h00050413,
32'h00044503,
32'h00051a63,
32'h00813083,
32'h00013403,
32'h01010113,
32'h00008067,
32'hfb9ff0ef,
32'h00140413,
32'hfe1ff06f,
32'hff010113,
32'h00113423,
32'hfc5ff0ef,
32'h00d00513,
32'hf9dff0ef,
32'h00813083,
32'h00a00513,
32'h01010113,
32'hf8dff06f,
32'hfd010113,
32'h02113423,
32'h00c13423,
32'h100247b7,
32'h00200713,
32'h02813023,
32'h00913c23,
32'h00e7ac23,
32'h00058413,
32'h00050493,
32'hf39ff0ef,
32'h00048513,
32'hf15ff0ef,
32'h0184551b,
32'hf0dff0ef,
32'h00000513,
32'hf05ff0ef,
32'h0084551b,
32'h0ff57513,
32'hef9ff0ef,
32'h0ff47513,
32'hef1ff0ef,
32'h00813503,
32'h3e800413,
32'hee5ff0ef,
32'hefdff0ef,
32'h0185179b,
32'h4187d79b,
32'h00050493,
32'h0007dc63,
32'hfff40413,
32'hfe0414e3,
32'h00000517,
32'h02c50513,
32'hf55ff0ef,
32'h02813083,
32'h02013403,
32'h00048513,
32'h01813483,
32'h03010113,
32'h00008067,
32'hf39ff06f,
32'h00000000,
32'h635f6473,
32'h203a646d,
32'h656d6974,
32'h0074756f,
32'h54494e49,
32'h00000000,
32'h00000000,
32'h00000000,
32'h30444d43,
32'h00000000,
32'h38444d43,
32'h00000000,
32'h444d4341,
32'h00003134,
32'h35444d43,
32'h00000038,
32'h31444d43,
32'h00000036,
32'h31444d43,
32'h00000038,
32'h44414f4c,
32'h20474e49,
32'h00000020,
32'h00000000,
32'h43202d08,
32'h6d204352,
32'h616d7369,
32'h20686374,
32'h00000000,
32'h00000000,
32'h00002008,
32'h00000000,
32'h4f525245,
32'h00000052,
32'h544f4f42


    };
    always_ff @(posedge clk or negedge rstn)
        if (!rstn)
            rvalid <= 1'b0;
        else
            rvalid <= addr_valid & addr_ready;

    always_ff @(posedge clk or negedge rstn)
        if (!rstn)
            rdata <= '0;
        else if (addr_valid & addr_ready)
            rdata <= rom_content[addr[31:2]];
    always_ff @(posedge clk or negedge rstn)
        if (!rstn)
            rdata2 <= '0;
        else if (addr2_valid & addr2_ready)
            rdata2 <= {rom_content[{addr2[31:3], 1'b1}], rom_content[{addr2[31:3], 1'b0}]};
    always_ff @(posedge clk or negedge rstn)
        if (!rstn)
            rvalid2 <= 1'b0;
        else
            rvalid2 <= addr2_valid & addr2_ready;
    assign addr_ready = 1'b1;
    assign addr2_ready = 1'b1;

endmodule